module skullart (vssd1, vccd1);
 input vssd1;
 input vccd1;
endmodule

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullart
  CLASS BLOCK ;
  FOREIGN skullart ;
  ORIGIN -10.000 -10.000 ;
  SIZE 90.000 BY 125.700 ;
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 95.000 10.000 100.000 135.700 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 10.000 10.000 15.000 135.700 ;
    END
  END vccd1
  OBS
      LAYER met1 ;
        RECT 47.300 133.000 68.900 135.700 ;
        RECT 44.600 130.300 68.900 133.000 ;
        RECT 39.200 124.900 74.300 130.300 ;
        RECT 36.500 114.100 77.000 124.900 ;
        RECT 36.500 111.400 44.600 114.100 ;
        RECT 36.500 108.700 41.900 111.400 ;
        RECT 39.200 106.000 41.900 108.700 ;
        RECT 52.700 106.000 60.800 114.100 ;
        RECT 68.900 111.400 77.000 114.100 ;
        RECT 71.600 108.700 77.000 111.400 ;
        RECT 71.600 106.000 74.300 108.700 ;
        RECT 39.200 103.300 44.600 106.000 ;
        RECT 50.000 103.300 63.500 106.000 ;
        RECT 68.900 103.300 74.300 106.000 ;
        RECT 39.200 100.600 55.400 103.300 ;
        RECT 58.100 100.600 71.600 103.300 ;
        RECT 44.600 97.900 52.700 100.600 ;
        RECT 60.800 97.900 71.600 100.600 ;
        RECT 47.300 92.500 66.200 97.900 ;
        RECT 31.100 89.800 39.200 92.500 ;
        RECT 47.300 89.800 50.000 92.500 ;
        RECT 52.700 89.800 55.400 92.500 ;
        RECT 58.100 89.800 60.800 92.500 ;
        RECT 63.500 89.800 66.200 92.500 ;
        RECT 74.300 89.800 82.400 92.500 ;
        RECT 28.400 84.400 41.900 89.800 ;
        RECT 71.600 84.400 85.100 89.800 ;
        RECT 31.100 81.700 47.300 84.400 ;
        RECT 66.200 81.700 82.400 84.400 ;
        RECT 39.200 79.000 50.000 81.700 ;
        RECT 63.500 79.000 74.300 81.700 ;
        RECT 44.600 76.300 55.400 79.000 ;
        RECT 58.100 76.300 68.900 79.000 ;
        RECT 50.000 70.900 63.500 76.300 ;
        RECT 44.600 68.200 55.400 70.900 ;
        RECT 58.100 68.200 68.900 70.900 ;
        RECT 31.100 65.500 50.000 68.200 ;
        RECT 63.500 65.500 85.100 68.200 ;
        RECT 28.400 62.800 44.600 65.500 ;
        RECT 68.900 62.800 85.100 65.500 ;
        RECT 28.400 60.100 39.200 62.800 ;
        RECT 74.300 60.100 85.100 62.800 ;
        RECT 28.400 57.400 36.500 60.100 ;
        RECT 77.000 57.400 85.100 60.100 ;
        RECT 31.100 54.700 33.800 57.400 ;
        RECT 47.300 54.700 50.000 57.400 ;
        RECT 52.700 54.700 55.400 57.400 ;
        RECT 58.100 54.700 60.800 57.400 ;
        RECT 63.500 54.700 66.200 57.400 ;
        RECT 79.700 54.700 82.400 57.400 ;
        RECT 47.300 49.300 66.200 54.700 ;
        RECT 44.600 46.600 52.700 49.300 ;
        RECT 60.800 46.600 71.600 49.300 ;
        RECT 39.200 43.900 55.400 46.600 ;
        RECT 58.100 43.900 71.600 46.600 ;
        RECT 39.200 41.200 44.600 43.900 ;
        RECT 50.000 41.200 63.500 43.900 ;
        RECT 68.900 41.200 74.300 43.900 ;
        RECT 39.200 38.500 41.900 41.200 ;
        RECT 36.500 35.800 41.900 38.500 ;
        RECT 36.500 33.100 44.600 35.800 ;
        RECT 52.700 33.100 60.800 41.200 ;
        RECT 71.600 38.500 74.300 41.200 ;
        RECT 71.600 35.800 77.000 38.500 ;
        RECT 68.900 33.100 77.000 35.800 ;
        RECT 36.500 22.300 77.000 33.100 ;
        RECT 39.200 16.900 74.300 22.300 ;
        RECT 44.600 14.200 68.900 16.900 ;
        RECT 47.300 11.500 68.900 14.200 ;
      LAYER met4 ;
        RECT 47.300 133.000 68.900 135.700 ;
        RECT 44.600 130.300 68.900 133.000 ;
        RECT 39.200 124.900 74.300 130.300 ;
        RECT 36.500 114.100 77.000 124.900 ;
        RECT 36.500 111.400 44.600 114.100 ;
        RECT 36.500 108.700 41.900 111.400 ;
        RECT 39.200 106.000 41.900 108.700 ;
        RECT 52.700 106.000 60.800 114.100 ;
        RECT 68.900 111.400 77.000 114.100 ;
        RECT 71.600 108.700 77.000 111.400 ;
        RECT 71.600 106.000 74.300 108.700 ;
        RECT 39.200 103.300 44.600 106.000 ;
        RECT 50.000 103.300 63.500 106.000 ;
        RECT 68.900 103.300 74.300 106.000 ;
        RECT 39.200 100.600 55.400 103.300 ;
        RECT 58.100 100.600 71.600 103.300 ;
        RECT 44.600 97.900 52.700 100.600 ;
        RECT 60.800 97.900 71.600 100.600 ;
        RECT 47.300 92.500 66.200 97.900 ;
        RECT 31.100 89.800 39.200 92.500 ;
        RECT 47.300 89.800 50.000 92.500 ;
        RECT 52.700 89.800 55.400 92.500 ;
        RECT 58.100 89.800 60.800 92.500 ;
        RECT 63.500 89.800 66.200 92.500 ;
        RECT 74.300 89.800 82.400 92.500 ;
        RECT 28.400 84.400 41.900 89.800 ;
        RECT 71.600 84.400 85.100 89.800 ;
        RECT 31.100 81.700 47.300 84.400 ;
        RECT 66.200 81.700 82.400 84.400 ;
        RECT 39.200 79.000 50.000 81.700 ;
        RECT 63.500 79.000 74.300 81.700 ;
        RECT 44.600 76.300 55.400 79.000 ;
        RECT 58.100 76.300 68.900 79.000 ;
        RECT 50.000 70.900 63.500 76.300 ;
        RECT 44.600 68.200 55.400 70.900 ;
        RECT 58.100 68.200 68.900 70.900 ;
        RECT 31.100 65.500 50.000 68.200 ;
        RECT 63.500 65.500 85.100 68.200 ;
        RECT 28.400 62.800 44.600 65.500 ;
        RECT 68.900 62.800 85.100 65.500 ;
        RECT 28.400 60.100 39.200 62.800 ;
        RECT 74.300 60.100 85.100 62.800 ;
        RECT 28.400 57.400 36.500 60.100 ;
        RECT 77.000 57.400 85.100 60.100 ;
        RECT 31.100 54.700 33.800 57.400 ;
        RECT 47.300 54.700 50.000 57.400 ;
        RECT 52.700 54.700 55.400 57.400 ;
        RECT 58.100 54.700 60.800 57.400 ;
        RECT 63.500 54.700 66.200 57.400 ;
        RECT 79.700 54.700 82.400 57.400 ;
        RECT 47.300 49.300 66.200 54.700 ;
        RECT 44.600 46.600 52.700 49.300 ;
        RECT 60.800 46.600 71.600 49.300 ;
        RECT 39.200 43.900 55.400 46.600 ;
        RECT 58.100 43.900 71.600 46.600 ;
        RECT 39.200 41.200 44.600 43.900 ;
        RECT 50.000 41.200 63.500 43.900 ;
        RECT 68.900 41.200 74.300 43.900 ;
        RECT 39.200 38.500 41.900 41.200 ;
        RECT 36.500 35.800 41.900 38.500 ;
        RECT 36.500 33.100 44.600 35.800 ;
        RECT 52.700 33.100 60.800 41.200 ;
        RECT 71.600 38.500 74.300 41.200 ;
        RECT 71.600 35.800 77.000 38.500 ;
        RECT 68.900 33.100 77.000 35.800 ;
        RECT 36.500 22.300 77.000 33.100 ;
        RECT 39.200 16.900 74.300 22.300 ;
        RECT 44.600 14.200 68.900 16.900 ;
        RECT 47.300 11.500 68.900 14.200 ;
  END
END skullart
END LIBRARY

